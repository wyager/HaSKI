// Automatically generated Verilog-2001
module Hardware_ram_11(eta_i1
                      ,// clock
                      system1000
                      ,// asynchronous reset: active low
                      system1000_rstn
                      ,bodyVar_o);
  input [95:0] eta_i1;
  input system1000;
  input system1000_rstn;
  output [65:0] bodyVar_o;
  wire [0:0] x_0;
  wire [0:0] x_1;
  wire [63:0] bodyVar_2;
  wire [0:0] a8_3;
  wire [0:0] a7_4;
  wire signed [31:0] bodyVar_5;
  wire [0:0] bodyVar_6;
  wire [63:0] repANF_7;
  wire signed [31:0] wild_8;
  wire [0:0] x_9;
  wire [0:0] x_10;
  wire [0:0] x_11;
  wire [0:0] x_12;
  wire signed [31:0] repANF_13;
  wire [63:0] x_14;
  wire [29:0] a9_15;
  wire [29:0] x_16;
  wire [0:0] tmp_17;
  wire [0:0] tmp_21;
  wire [63:0] tmp_25;
  wire signed [31:0] tmp_72;
  assign bodyVar_o = {x_0
                     ,x_1
                     ,bodyVar_2};
  
  // register begin
  reg [0:0] n_19;
  
  always @(posedge system1000 or negedge system1000_rstn) begin : register_Hardware_ram_11_n_20
    if (~ system1000_rstn) begin
      n_19 <= 1'b0;
    end else begin
      n_19 <= a7_4;
    end
  end
  
  assign tmp_17 = n_19;
  // register end
  
  assign x_0 = tmp_17;
  
  // register begin
  reg [0:0] n_23;
  
  always @(posedge system1000 or negedge system1000_rstn) begin : register_Hardware_ram_11_n_24
    if (~ system1000_rstn) begin
      n_23 <= 1'b0;
    end else begin
      n_23 <= a8_3;
    end
  end
  
  assign tmp_21 = n_23;
  // register end
  
  assign x_1 = tmp_21;
  
  // blockRam begin
  reg [63:0] RAM_n_65 [0:1280-1];
  reg [63:0] dout_n_66;
  
  reg [81919:0] ram_init_n_67;
  integer n_68;
  initial begin
    ram_init_n_67 = ({{64'b0011000000000000000000000000000001000000000000000000000000000110,64'b0011000000000000000000000000000010000000000000000000000000000101,64'b0011000000000000000000000000000011000000000000000000000000000100,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0010000000000000000000000000000000000000000000000000000000000000,64'b0010000000000000000000000000000000000000000000000000000000000000,64'b0011000000000000000000000000000111000000000000000000000000001100,64'b0011000000000000000000000000001000000000000000000000000000001011,64'b0011000000000000000000000000001001000000000000000000000000001010,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0010000000000000000000000000000000000000000000000000000000000000,64'b0010000000000000000000000000000000000000000000000000000000000000,64'b0011000000000000000000000000001101000000000000000000000000100010,64'b0011000000000000000000000000001110000000000000000000000000100001,64'b0011000000000000000000000000001111000000000000000000000000100000,64'b0011000000000000000000000000010000000000000000000000000000011111,64'b0011000000000000000000000000010001000000000000000000000000011110,64'b0011000000000000000000000000010010000000000000000000000000011101,64'b0011000000000000000000000000010011000000000000000000000000011100,64'b0011000000000000000000000000010100000000000000000000000000011011,64'b0011000000000000000000000000010101000000000000000000000000011010,64'b0011000000000000000000000000010110000000000000000000000000011001,64'b0011000000000000000000000000010111000000000000000000000000011000,64'b0100000000000000000000000000000000000000000000000000000001101000,64'b0100000000000000000000000000000000000000000000000000000001100101,64'b0100000000000000000000000000000000000000000000000000000001101100,64'b0100000000000000000000000000000000000000000000000000000001101100,64'b0100000000000000000000000000000000000000000000000000000001101111,64'b0100000000000000000000000000000000000000000000000000000001011111,64'b0100000000000000000000000000000000000000000000000000000001110111,64'b0100000000000000000000000000000000000000000000000000000001101111,64'b0100000000000000000000000000000000000000000000000000000001110010,64'b0100000000000000000000000000000000000000000000000000000001101100,64'b0100000000000000000000000000000000000000000000000000000001100100,64'b0100000000000000000000000000000000000000000000000000000000100001},({(1245) {64'b0000000000000000000000000000000000000000000000000000000000000000}})});
    for (n_68=0; n_68 < 1280; n_68 = n_68 + 1) begin
      RAM_n_65[1280-1-n_68] = ram_init_n_67[n_68*64+:64];
    end
  end
  
  always @(posedge system1000) begin : blockRam_Hardware_ram_11_n_69
    if (bodyVar_6) begin
      RAM_n_65[bodyVar_5] <= repANF_7;
    end
    dout_n_66 <= RAM_n_65[bodyVar_5];
  end
  
  assign tmp_25 = dout_n_66;
  // blockRam end
  
  assign bodyVar_2 = tmp_25;
  
  assign a8_3 = x_11;
  
  assign a7_4 = x_12;
  
  assign bodyVar_5 = wild_8;
  
  assign bodyVar_6 = x_9 & x_10;
  
  assign repANF_7 = x_14;
  
  assign wild_8 = repANF_13;
  
  Hardware_ram1_12 Hardware_ram1_12_x_9
  (.topLet_o (x_9)
  ,.ds1_i1 (a7_4));
  
  Hardware_ram1_12 Hardware_ram1_12_x_10
  (.topLet_o (x_10)
  ,.ds1_i1 (a8_3));
  
  assign x_11 = eta_i1[94:94];
  
  assign x_12 = eta_i1[95:95];
  
  assign tmp_72 = $unsigned(a9_15);
  
  assign repANF_13 = tmp_72;
  
  assign x_14 = eta_i1[63:0];
  
  assign a9_15 = x_16;
  
  assign x_16 = eta_i1[93:64];
endmodule
