// Automatically generated Verilog-2001
module Hardware_topEntity(// clock
                         system1000
                         ,// asynchronous reset: active low
                         system1000_rstn
                         ,output_0_0_0
                         ,output_0_0_1
                         ,output_0_1);
  input system1000;
  input system1000_rstn;
  output [0:0] output_0_0_0;
  output [31:0] output_0_0_1;
  output [0:0] output_0_1;
  wire [33:0] output_0;
  wire [32:0] output_0_0;
  Hardware_topEntity_0 Hardware_topEntity_0_inst
  (.system1000 (system1000)
  ,.system1000_rstn (system1000_rstn)
  ,.topLet_o (output_0));
  
  assign output_0_0 = output_0[33:1];
  
  assign output_0_1 = output_0[0:0];
  
  assign output_0_0_0 = output_0_0[32:32];
  
  assign output_0_0_1 = output_0_0[31:0];
endmodule
