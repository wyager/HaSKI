// Automatically generated Verilog-2001
module Hardware_ram_11(eta_i1
                      ,// clock
                      system1000
                      ,// asynchronous reset: active low
                      system1000_rstn
                      ,y_o);
  input [95:0] eta_i1;
  input system1000;
  input system1000_rstn;
  output [65:0] y_o;
  wire [32833:0] altLet_0;
  wire [95:0] x_1;
  wire [32833:0] bodyVar_2;
  wire [32833:0] altLet_3;
  wire [0:0] ds2_4;
  wire [95:0] repANF_5;
  wire [32833:0] altLet_6;
  wire [32767:0] x_7;
  wire [32833:0] altLet_8;
  wire [32833:0] altLet_9;
  wire [0:0] ds3_10;
  wire [65:0] repANF_11;
  wire [32767:0] bodyVar_12;
  wire [63:0] bodyVar_13;
  wire [63:0] ds5_14;
  wire [32767:0] x_15;
  wire signed [31:0] repANF_16;
  wire signed [31:0] wild5_17;
  wire signed [31:0] repANF_18;
  wire [29:0] ds4_19;
  wire [95:0] tmp_20;
  wire [95:0] tmp_31;
  wire [32767:0] tmp_39;
  wire [32767:0] tmp_86;
  wire [63:0] tmp_92;
  wire signed [31:0] tmp_98;
  assign y_o = altLet_0[65:0];
  
  reg [32833:0] altLet_0_reg;
  always @(*) begin
    case(ds2_4)
      1'b0 : altLet_0_reg = altLet_3;
      default : altLet_0_reg = bodyVar_2;
    endcase
  end
  assign altLet_0 = altLet_0_reg;
  
  // register begin
  reg [95:0] n_25;
  
  always @(posedge system1000 or negedge system1000_rstn) begin : register_Hardware_ram_11_n_26
    if (~ system1000_rstn) begin
      n_25 <= {1'b0,1'b0,30'b000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
    end else begin
      n_25 <= repANF_5;
    end
  end
  
  assign tmp_20 = n_25;
  // register end
  
  assign x_1 = tmp_20;
  
  reg [32833:0] bodyVar_2_reg;
  always @(*) begin
    case(ds2_4)
      1'b1 : bodyVar_2_reg = altLet_6;
      default : bodyVar_2_reg = {32834 {1'bx}};
    endcase
  end
  assign bodyVar_2 = bodyVar_2_reg;
  
  assign altLet_3 = {x_7
                    ,{1'b0
                     ,1'b0
                     ,64'b0000000000000000000000000000000000000000000000000000000000000000}};
  
  assign ds2_4 = x_1[95:95];
  
  // register begin
  reg [95:0] n_36;
  
  always @(posedge system1000 or negedge system1000_rstn) begin : register_Hardware_ram_11_n_37
    if (~ system1000_rstn) begin
      n_36 <= {1'b0,1'b0,30'b000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
    end else begin
      n_36 <= eta_i1;
    end
  end
  
  assign tmp_31 = n_36;
  // register end
  
  assign repANF_5 = tmp_31;
  
  reg [32833:0] altLet_6_reg;
  always @(*) begin
    case(ds3_10)
      1'b0 : altLet_6_reg = altLet_8;
      1'b1 : altLet_6_reg = altLet_9;
      default : altLet_6_reg = {32834 {1'bx}};
    endcase
  end
  assign altLet_6 = altLet_6_reg;
  
  // register begin
  reg [32767:0] n_79;
  
  always @(posedge system1000 or negedge system1000_rstn) begin : register_Hardware_ram_11_n_80
    if (~ system1000_rstn) begin
      n_79 <= ({{64'b0011000000000000000000000000000001000000000000000000000000000110,64'b0011000000000000000000000000000010000000000000000000000000000101,64'b0011000000000000000000000000000011000000000000000000000000000100,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0010000000000000000000000000000000000000000000000000000000000000,64'b0010000000000000000000000000000000000000000000000000000000000000,64'b0011000000000000000000000000000111000000000000000000000000001100,64'b0011000000000000000000000000001000000000000000000000000000001011,64'b0011000000000000000000000000001001000000000000000000000000001010,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0010000000000000000000000000000000000000000000000000000000000000,64'b0010000000000000000000000000000000000000000000000000000000000000,64'b0011000000000000000000000000001101000000000000000000000000100010,64'b0011000000000000000000000000001110000000000000000000000000100001,64'b0011000000000000000000000000001111000000000000000000000000100000,64'b0011000000000000000000000000010000000000000000000000000000011111,64'b0011000000000000000000000000010001000000000000000000000000011110,64'b0011000000000000000000000000010010000000000000000000000000011101,64'b0011000000000000000000000000010011000000000000000000000000011100,64'b0011000000000000000000000000010100000000000000000000000000011011,64'b0011000000000000000000000000010101000000000000000000000000011010,64'b0011000000000000000000000000010110000000000000000000000000011001,64'b0011000000000000000000000000010111000000000000000000000000011000,64'b0100000000000000000000000000000000000000000000000000000001101000,64'b0100000000000000000000000000000000000000000000000000000001100101,64'b0100000000000000000000000000000000000000000000000000000001101100,64'b0100000000000000000000000000000000000000000000000000000001101100,64'b0100000000000000000000000000000000000000000000000000000001101111,64'b0100000000000000000000000000000000000000000000000000000001011111,64'b0100000000000000000000000000000000000000000000000000000001110111,64'b0100000000000000000000000000000000000000000000000000000001101111,64'b0100000000000000000000000000000000000000000000000000000001110010,64'b0100000000000000000000000000000000000000000000000000000001101100,64'b0100000000000000000000000000000000000000000000000000000001100100,64'b0100000000000000000000000000000000000000000000000000000000100001},({(477) {64'b0000000000000000000000000000000000000000000000000000000000000000}})});
    end else begin
      n_79 <= x_15;
    end
  end
  
  assign tmp_39 = n_79;
  // register end
  
  assign x_7 = tmp_39;
  
  assign altLet_8 = {x_7
                    ,repANF_11};
  
  assign altLet_9 = {bodyVar_12
                    ,{1'b1
                     ,1'b1
                     ,64'b0000000000000000000000000000000000000000000000000000000000000000}};
  
  assign ds3_10 = x_1[94:94];
  
  assign repANF_11 = {1'b1
                     ,1'b0
                     ,bodyVar_13};
  
  // replaceVec start
  wire [32767:0] vecflat_n_87;
  assign vecflat_n_87 = x_7;
  
  reg [63:0] vec_n_88 [0:512-1];
  integer n_89;
  always @(*) begin
    for (n_89=0;n_89<512;n_89=n_89+1) begin
      vec_n_88[512-1-n_89] = vecflat_n_87[n_89*64+:64];
    end
    vec_n_88[repANF_16] = ds5_14;
  end
  
  genvar n_90;
  generate
  for (n_90=0;n_90<512;n_90=n_90+1) begin : vec_n_91
    assign tmp_86[n_90*64+:64] = vec_n_88[(512-1)-n_90];
  end
  endgenerate
  // replaceVec end
  
  assign bodyVar_12 = tmp_86;
  
  // indexVec begin
  wire [63:0] vec_n_93 [0:512-1];
  
  wire [32767:0] vecflat_n_94;
  assign vecflat_n_94 = x_7;
  genvar n_95;
  generate
  for (n_95=0; n_95 < 512; n_95=n_95+1) begin : array_n_96
    assign vec_n_93[(512-1)-n_95] = vecflat_n_94[n_95*64+:64];
  end
  endgenerate
  
  assign tmp_92 = vec_n_93[repANF_16];
  // indexVec end
  
  assign bodyVar_13 = tmp_92;
  
  assign ds5_14 = x_1[63:0];
  
  assign x_15 = altLet_0[32833:66];
  
  assign repANF_16 = wild5_17;
  
  assign wild5_17 = repANF_18;
  
  assign tmp_98 = $unsigned(ds4_19);
  
  assign repANF_18 = tmp_98;
  
  assign ds4_19 = x_1[93:64];
endmodule
