// Automatically generated Verilog-2001
module Hardware_topEntity_0(// clock
                           system1000
                           ,// asynchronous reset: active low
                           system1000_rstn
                           ,topLet_o);
  input system1000;
  input system1000_rstn;
  output [33:0] topLet_o;
  wire [32:0] repANF_0;
  wire [0:0] repANF_1;
  Hardware_topEntity7_1 Hardware_topEntity7_1_repANF_0
  (.topLet_o (repANF_0)
  ,.system1000 (system1000)
  ,.system1000_rstn (system1000_rstn));
  
  Hardware_topEntity1_15 Hardware_topEntity1_15_repANF_1
  (.topLet_o (repANF_1)
  ,.system1000 (system1000)
  ,.system1000_rstn (system1000_rstn));
  
  assign topLet_o = {repANF_0
                    ,repANF_1};
endmodule
